library verilog;
use verilog.vl_types.all;
entity CentralProcessorUnit is
end CentralProcessorUnit;
