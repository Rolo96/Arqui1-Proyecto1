library verilog;
use verilog.vl_types.all;
entity CentralProcessorUnit_tb is
end CentralProcessorUnit_tb;
