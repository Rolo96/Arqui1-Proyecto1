`timescale 1ns / 1ps
module CentralProcessorUnit();

endmodule
