`timescale 1ns / 1ps
module CentralProcessorUnit_tb();

endmodule